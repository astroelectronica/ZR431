.title KiCad schematic
.include "C:/AE/ZR431/_models/BAS21.spice.txt"
.include "C:/AE/ZR431/_models/C1608C0G1H470J080AA_p.mod"
.include "C:/AE/ZR431/_models/C2012X5R1E106M125AB_p.mod"
.include "C:/AE/ZR431/_models/FMMT493.spice.txt"
.include "C:/AE/ZR431/_models/ZR431.spice.txt"
XU3 /VOUT 0 C2012X5R1E106M125AB_p
I1 /VOUT 0 {ILOAD}
R1 /VC /VZ {RBASE}
V1 /VIN 0 {VSOURCE}
D1 /VIN /VC DI_BAS21
XU1 /VZ /VREF C1608C0G1H470J080AA_p
R3 /VREF 0 {RREF}
R2 /VOUT /VREF {RADJ}
Q1 /VC /VZ /VOUT FMMT493
XU2 /VZ /VREF 0 ZR431
.end
